package data_types is
  type stav_t is (RES,STARTING,WAITING,STORE,COMP,PUSH);
end data_types;
