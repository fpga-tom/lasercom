package data_types is
  type stav_t is (RES,STARTING,LOAD,STORE,COMP,PUSH);
end data_types;
